-------------------------------------------------------------------------
-- Henry Duwe
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------
-- MIPS_Processor.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a skeleton of a MIPS_Processor  
-- implementation.
-- 01/29/2019 by H3::Design created.
-------------------------------------------------------------------------

library IEEE;
  use IEEE.std_logic_1164.all;

library work;
  use work.MIPS_types.all;

entity MIPS_Processor is
  generic (N : integer := DATA_WIDTH);
  port (iCLK      : in  std_logic;
        iRST      : in  std_logic;
        iInstLd   : in  std_logic;
        iInstAddr : in  std_logic_vector(N - 1 downto 0);
        iInstExt  : in  std_logic_vector(N - 1 downto 0);
        oALUOut   : out std_logic_vector(N - 1 downto 0)); -- TODO: Hook this up to the output of the ALU. It is important for synthesis that you have this output that can effectively be impacted by all other components so they are not optimized away.

end entity;

architecture structure of MIPS_Processor is

  component mem is
    generic (ADDR_WIDTH : integer;
             DATA_WIDTH : integer);
    port (
      clk  : in  std_logic;
      addr : in  std_logic_vector((ADDR_WIDTH - 1) downto 0);
      data : in  std_logic_vector((DATA_WIDTH - 1) downto 0);
      we   : in  std_logic := '1';
      q    : out std_logic_vector((DATA_WIDTH - 1) downto 0));
  end component;

  component ALU is
    port (i_ALU_A        : in  std_logic_vector(N - 1 downto 0); -- ALU Input A
          i_ALU_B        : in  std_logic_vector(N - 1 downto 0); -- ALU Input B
          i_ALU_Ctl      : in  std_logic_vector(4 downto 0);     -- ALU Control Input [4]Signed or unsidned, [3]shift L or A, [2]selector, [1]selector, [0]selector
          o_ALU_Carry    : out std_logic;                        -- ALU Indicator for a carry out bit.
          o_ALU_Zero     : out std_logic;                        -- ALU Indicator that an operation has resulting in a 0 output.
          o_ALU_Overflow : out std_logic;                        -- ALU Indicator that an overflow has occured.
          o_ALU_I_Result : out std_logic_vector(N - 1 downto 0)); -- ALU add Sub Results.
  end component;

  component AdderSubtractor is
    port (i_AddSub_A        : in  std_logic_vector(N - 1 downto 0);
          i_AddSub_B        : in  std_logic_vector(N - 1 downto 0);
          i_AddSub_nAdd_sub : in  std_logic;
          o_AddSub_Sum      : out std_logic_vector(N - 1 downto 0);
          o_AddSub_Cout     : out std_logic;
          o_AddSub_Overflow : out std_logic;
          o_AddSub_Zero     : out std_logic);
  end component;

  component RippleCarryAdder is
    port (A        : in  std_logic_vector(N - 1 downto 0);
          B        : in  std_logic_vector(N - 1 downto 0);
          Sum      : out std_logic_vector(N - 1 downto 0);
          Carry    : out std_logic; -- Final carry out
          --           Zero    : out std_logic; -- Indicates if Sum is zero
          Overflow : out std_logic); -- Indicates overflow condition
  end component;

  component OnesComplementor is
    port (i_D0 : in  std_logic_vector(N - 1 downto 0);
          o_O  : out std_logic_vector(N - 1 downto 0));
  end component;

  component Shifter is
    port (i_in        : in  std_logic_vector(N - 1 downto 0);
          i_shift_C   : in  std_logic; --0 = Logical, 1 = Arithmetic
          i_Direction : in  std_logic; --0 = left, 1 = right
          i_Shamt     : in  std_logic_vector(4 downto 0);
          o_Out       : out std_logic_vector(N - 1 downto 0));
  end component;

  component mux2t1_N is
    port (
      i_s  : in  std_logic;
      i_D0 : in  std_logic_vector(N - 1 downto 0);
      i_D1 : in  std_logic_vector(N - 1 downto 0);
      o_O  : out std_logic_vector(N - 1 downto 0)
    );
  end component;

  component mux8t1_N is
    port (i_w0, i_w1, i_w2, i_w3 : in  std_logic_vector(N - 1 downto 0);
          i_w4, i_w5, i_w6, i_w7 : in  std_logic_vector(N - 1 downto 0);
          i_s0                   : in  std_logic;
          i_s1                   : in  std_logic;
          i_s2                   : in  std_logic;
          o_Y                    : out std_logic_vector(N - 1 downto 0));
  end component;

  component fetchLogic is
    port (
      i_jump_C          : in  std_logic;
      i_jr_ra_C         : in  std_logic;
      i_CLK             : in  std_logic;
      i_RST             : in  std_logic;
      i_w_branch_n_ALUo : in  std_logic;
      i_instr_25t0      : in  std_logic_vector(25 downto 0);
      i_ext_imm         : in  std_logic_vector(N - 1 downto 0);
      i_jr_ra_pc_next   : in  std_logic_vector(N - 1 downto 0);
      o_pc_p4           : out std_logic_vector(N - 1 downto 0);
      o_pc_next         : out std_logic_vector(N - 1 downto 0));
  end component;

  component controller is
    port (i_instruct31_26 : in  std_logic_vector(5 downto 0);
          i_instruct5_0   : in  std_logic_vector(5 downto 0);
          o_STD_SHIFT     : out std_logic; -- Standard shift (1)we are doing a normal shift (0) we are doing a variable shift or does not matter.
          o_ALU_Ctl       : out std_logic_vector(4 downto 0);
          o_RegWrite      : out std_logic;
          o_MemtoReg      : out std_logic;
          o_MemWrite      : out std_logic;
          o_MemRead       : out std_logic;
          o_RegDst        : out std_logic_vector(1 downto 0);
          o_Branch        : out std_logic;
          o_Alu_Src       : out std_logic;
          o_ext_ctl       : out std_logic;
          o_Jump          : out std_logic;
          o_jr            : out std_logic;
          o_jal           : out std_logic);
  end component;

  -- Required data memory signals
  signal s_DMemWr   : std_logic;                        -- TODO: use this signal as the final active high data memory write enable signal
  signal s_DMemAddr : std_logic_vector(N - 1 downto 0); -- TODO: use this signal as the final data memory address input
  signal s_DMemData : std_logic_vector(N - 1 downto 0); -- TODO: use this signal as the final data memory data input
  signal s_DMemOut  : std_logic_vector(N - 1 downto 0); -- TODO: use this signal as the data memory output

  -- Required register file signals 
  signal s_RegWr     : std_logic;                        -- TODO: use this signal as the final active high write enable input to the register file
  signal s_RegWrAddr : std_logic_vector(4 downto 0);     -- TODO: use this signal as the final destination register address input
  signal s_RegWrData : std_logic_vector(N - 1 downto 0); -- TODO: use this signal as the final data memory data input

  -- Required instruction memory signals
  signal s_IMemAddr     : std_logic_vector(N - 1 downto 0); -- Do not assign this signal, assign to s_NextInstAddr instead
  signal s_NextInstAddr : std_logic_vector(N - 1 downto 0); -- TODO: use this signal as your intended final instruction memory address input.
  signal s_Inst         : std_logic_vector(N - 1 downto 0); -- TODO: use this signal as the instruction signal 

  -- Required halt signal -- for simulation
  signal s_Halt : std_logic; -- TODO: this signal indicates to the simulation that intended program execution has completed. (Opcode: 01 0100)

  -- Required overflow signal -- for overflow exception detection
  signal s_Ovfl : std_logic; -- TODO: this signal indicates an overflow exception would have been initiated

  -- TODO: You may add any additional signals or components your implementation 
  --       requires below this comment

begin

  -- TODO: This is required to be your final input to your instruction memory. This provides a feasible method to externally load the memory module which means that the synthesis tool must assume it knows nothing about the values stored in the instruction memory. If this is not included, much, if not all of the design is optimized out because the synthesis tool will believe the memory to be all zeros.
  with iInstLd select
    s_IMemAddr <= s_NextInstAddr when '0',
                  iInstAddr      when others;

  IMem: mem
    generic map (ADDR_WIDTH => ADDR_WIDTH,
                 DATA_WIDTH => N)
    port map (clk  => iCLK,
              addr => s_IMemAddr(11 downto 2),
              data => iInstExt,
              we   => iInstLd,
              q    => s_Inst);

  DMem: mem
    generic map (ADDR_WIDTH => ADDR_WIDTH,
                 DATA_WIDTH => N)
    port map (clk  => iCLK,
              addr => s_DMemAddr(11 downto 2),
              data => s_DMemData,
              we   => s_DMemWr,
              q    => s_DMemOut);

  -- TODO: Ensure that s_Halt is connected to an output control signal produced from decoding the Halt instruction (Opcode: 01 0100)
  -- TODO: Ensure that s_Ovfl is connected to the overflow output of your ALU
  -- TODO: Implement the rest of your processor below this comment! 
end architecture;

